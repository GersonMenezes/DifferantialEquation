library verilog;
use verilog.vl_types.all;
entity Multiplicador_Matricial_vlg_vec_tst is
end Multiplicador_Matricial_vlg_vec_tst;
