library verilog;
use verilog.vl_types.all;
entity Multiplicador_Matricial_vlg_check_tst is
    port(
        s               : in     vl_logic_vector(15 downto 0);
        sampler_rx      : in     vl_logic
    );
end Multiplicador_Matricial_vlg_check_tst;
