library verilog;
use verilog.vl_types.all;
entity DifferentialEquation_vlg_vec_tst is
end DifferentialEquation_vlg_vec_tst;
